
module empty();

endmodule
