module simple_comb_neg(
  input i,
  output o
);

assign o = ~i;

endmodule
