module verinject_mem1_injector
#(parameter LEFT = 0, parameter RIGHT = 0,
  parameter ADDR_LEFT = 0, parameter ADDR_RIGHT = 0,
  parameter MEM_LEFT = 0, parameter MEM_RIGHT = 0,
  parameter P_START = 0)
(
  // injector parameters
  input [31:0] verinject__injector_state,
  // clocking
  input clock,
  // memory read injection
  input [LEFT:RIGHT] unmodified,
  input [ADDR_LEFT:ADDR_RIGHT] read_address,
  output reg [LEFT:RIGHT] modified,
  // memory write capture
  input do_write,
  input [ADDR_LEFT:ADDR_RIGHT] write_address
);

wire [31:0] bits_start;
assign bits_start = (LEFT < RIGHT) ? LEFT : RIGHT;
wire [31:0] word_len;
assign word_len = (LEFT < RIGHT) ? (RIGHT - LEFT + 1) : (LEFT - RIGHT + 1);
wire [31:0] mem_start;
assign mem_start = (MEM_LEFT < MEM_RIGHT) ? MEM_LEFT : MEM_RIGHT;
wire [31:0] mem_len;
assign mem_len = (MEM_LEFT < MEM_RIGHT) ? (MEM_RIGHT - MEM_LEFT + 1) : (MEM_LEFT - MEM_RIGHT + 1);

wire [31:0] read_word_start;
wire [31:0] read_word_end;
assign read_word_start = P_START + (read_address - mem_start) * word_len;
assign read_word_end = read_word_start + word_len;

reg [LEFT:RIGHT] xor_modifier;

always @*
begin : fault_injection
  modified = unmodified;
  if (verinject__injector_state >= read_word_start && verinject__injector_state < read_word_end)
  begin
    xor_modifier = (1 << (verinject__injector_state - read_word_start + bits_start));
    modified = unmodified ^ xor_modifier;
  end
end

endmodule
