
module empty(input a);

endmodule
